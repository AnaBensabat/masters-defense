<?xml version="1.0" encoding="UTF-8" standalone="no"?>
<!-- Created with Inkscape (http://www.inkscape.org/) -->

<svg
   width="179.22353mm"
   height="180.73051mm"
   viewBox="0 0 179.22353 180.73053"
   version="1.1"
   id="svg1"
   inkscape:version="1.4.2 (ebf0e940d0, 2025-05-08)"
   sodipodi:docname="slide-13.svg"
   inkscape:export-filename="../slide-13.png"
   inkscape:export-xdpi="96"
   inkscape:export-ydpi="96"
   xmlns:inkscape="http://www.inkscape.org/namespaces/inkscape"
   xmlns:sodipodi="http://sodipodi.sourceforge.net/DTD/sodipodi-0.dtd"
   xmlns:xlink="http://www.w3.org/1999/xlink"
   xmlns="http://www.w3.org/2000/svg"
   xmlns:svg="http://www.w3.org/2000/svg"
   xmlns:ns58="http://www.iki.fi/pav/software/textext/">
  <sodipodi:namedview
     id="namedview1"
     pagecolor="#ffffff"
     bordercolor="#000000"
     borderopacity="0.25"
     inkscape:showpageshadow="2"
     inkscape:pageopacity="0.0"
     inkscape:pagecheckerboard="0"
     inkscape:deskcolor="#d1d1d1"
     inkscape:document-units="mm"
     inkscape:zoom="0.66016601"
     inkscape:cx="78.010681"
     inkscape:cy="438.52606"
     inkscape:window-width="1876"
     inkscape:window-height="1006"
     inkscape:window-x="0"
     inkscape:window-y="0"
     inkscape:window-maximized="1"
     inkscape:current-layer="svg1">
    <inkscape:page
       x="0"
       y="0"
       width="179.22353"
       height="180.73053"
       id="page2"
       margin="0"
       bleed="0" />
  </sodipodi:namedview>
  <defs
     id="defs1">
    <marker
       style="overflow:visible"
       id="marker227"
       refX="0"
       refY="0"
       orient="auto"
       inkscape:stockid="Stop"
       markerWidth="0.64999998"
       markerHeight="0.64999998"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         style="fill:none;stroke:context-stroke;stroke-width:1"
         d="M 0,4 V -4"
         id="path227" />
    </marker>
    <marker
       style="overflow:visible"
       id="Stop"
       refX="0"
       refY="0"
       orient="auto"
       inkscape:stockid="Stop"
       markerWidth="0.64999998"
       markerHeight="0.64999998"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         style="fill:none;stroke:context-stroke;stroke-width:1"
         d="M 0,4 V -4"
         id="path23" />
    </marker>
    <inkscape:perspective
       sodipodi:type="inkscape:persp3d"
       inkscape:vp_x="-33.340517 : 9.3825959 : 0"
       inkscape:vp_y="0 : 318.01552 : 0"
       inkscape:vp_z="186.59184 : 66.406508 : 1"
       inkscape:persp3d-origin="153.25132 : 57.023914 : 1"
       id="perspective219" />
    <linearGradient
       id="linearGradient13"
       inkscape:collect="always">
      <stop
         style="stop-color:#9d552b;stop-opacity:0.96078431;"
         offset="0.92472827"
         id="stop13" />
      <stop
         style="stop-color:#9d552b;stop-opacity:0;"
         offset="1"
         id="stop14" />
    </linearGradient>
    <marker
       style="overflow:visible"
       id="marker13"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Wide arrow"
       markerWidth="1"
       markerHeight="1"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         style="fill:none;stroke:context-stroke;stroke-width:1;stroke-linecap:butt"
         d="M 3,-3 0,0 3,3"
         transform="rotate(180,0.125,0)"
         sodipodi:nodetypes="ccc"
         id="path13" />
    </marker>
    <marker
       style="overflow:visible"
       id="ArrowWide"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Wide arrow"
       markerWidth="1"
       markerHeight="1"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         style="fill:none;stroke:context-stroke;stroke-width:1;stroke-linecap:butt"
         d="M 3,-3 0,0 3,3"
         transform="rotate(180,0.125,0)"
         sodipodi:nodetypes="ccc"
         id="path12" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7" />
    </marker>
    <linearGradient
       id="linearGradient6"
       inkscape:collect="always">
      <stop
         style="stop-color:#000000;stop-opacity:1;"
         offset="0"
         id="stop6" />
      <stop
         style="stop-color:#000000;stop-opacity:0;"
         offset="1"
         id="stop7" />
    </linearGradient>
    <linearGradient
       id="linearGradient4"
       inkscape:collect="always">
      <stop
         style="stop-color:#0292b1;stop-opacity:0.58146107;"
         offset="0"
         id="stop3" />
      <stop
         style="stop-color:#004f59;stop-opacity:0.80780524;"
         offset="1"
         id="stop4" />
    </linearGradient>
    <linearGradient
       id="linearGradient1"
       inkscape:collect="always">
      <stop
         style="stop-color:#ea6502;stop-opacity:0.58146107;"
         offset="0"
         id="stop1" />
      <stop
         style="stop-color:#863100;stop-opacity:0.80780524;"
         offset="1"
         id="stop2" />
    </linearGradient>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient1"
       id="radialGradient2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="translate(-7.4238862,-2.4746288)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,27.481737,35.580308)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,34.218627,41.730806)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,27.835497,42.390374)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,40.146547,40.708026)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,36.439697,48.459854)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,36.262617,36.685338)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,10.186772,38.521799)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,23.019847,49.954473)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,14.431554,57.105742)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,44.007547,47.542068)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-8-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,42.798927,35.725655)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,64.26802,13.325055)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,67.53101,18.052198)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,8.1808838,76.069234)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,5.3058823,68.88318)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,48.943889,52.010858)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-1-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,49.623317,43.20815)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,40.641767,28.243798)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,51.174907,35.161077)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,30.742607,28.947029)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,20.242817,37.277741)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,21.568307,59.550384)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,36.387177,65.266406)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,50.36684,63.287898)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,22.843557,29.926935)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,58.170587,43.739513)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,24.350067,66.622308)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,16.128443,48.825108)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,17.690043,45.375014)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,53.520556,57.526792)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-24.301905,50.903016)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,13.213729,40.464467)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,16.629133,32.310385)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,32.653323,70.994156)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-69.455128,-32.912668)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-62.718238,-26.762168)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-38"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-76.694048,-31.215228)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,50.802731,-19.535464)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-47.744617,-16.083107)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,27.099822,27.576964)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-64"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-36.126298,-44.761146)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-36.363139,18.122676)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-04"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,64.237898,-63.64109)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-0-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-51.478471,-10.355357)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,20.890733,21.752214)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-1-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-66.194258,-39.545948)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-69.101368,-26.102598)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-56"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-73.917018,-18.538498)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,58.437973,-76.34595)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-52.176915,36.316774)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-49.397835,22.904835)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5-5-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,19.958441,-45.830826)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87-0-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,8.2244126,33.329116)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-8-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,22.837679,16.369144)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-8-6-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-42.768937,-3.6608305)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-5.1804232,-59.437171)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-1-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,28.824448,18.592674)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-1-3-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,20.615544,27.821274)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-60.674248,-31.807638)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-5-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-34.392957,-4.2254105)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-1-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-53.109579,64.839383)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-6-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-67.850318,-19.565678)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-79.246822,-23.117958)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-69.344375,60.029609)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-22.213367,52.296675)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-83.723136,-28.028508)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-8-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-80.307732,-36.182588)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-4-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,47.467667,67.077771)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,23.038779,53.277566)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,38.624584,67.596135)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,31.725155,50.350346)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,31.592641,49.615275)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-6-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,45.679543,53.852053)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-6-8-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,20.080548,61.719614)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.27800922,0,0,0.27800922,112.1701,-24.738724)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,30.583512,34.696294)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,41.636045,70.593289)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62-0-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,32.368976,10.494865)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62-0-9-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,67.179354,45.722457)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62-0-9-5-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,10.394666,35.036986)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-62-0-9-5-9-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,59.903104,46.175688)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-73.203144,57.924086)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-22.220241,64.435169)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-0-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-53.895848,14.9938)" />
    <linearGradient
       inkscape:collect="always"
       xlink:href="#linearGradient6"
       id="linearGradient7"
       x1="117.26712"
       y1="25.713768"
       x2="120.29007"
       y2="26.751619"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(2.733218,0,0,0.98185997,-190.32271,-43.697736)" />
    <marker
       style="overflow:visible"
       id="marker14-7"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Wide arrow"
       markerWidth="1"
       markerHeight="1"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         style="fill:none;stroke:context-stroke;stroke-width:1;stroke-linecap:butt"
         d="M 3,-3 0,0 3,3"
         transform="rotate(180,0.125,0)"
         sodipodi:nodetypes="ccc"
         id="path14-5" />
    </marker>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient13"
       id="radialGradient14"
       cx="43.384182"
       cy="44.199886"
       fx="43.384182"
       fy="44.199886"
       r="41.30278"
       gradientUnits="userSpaceOnUse" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-9-7"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.18455199,0,0,0.18455199,41.536591,-164.01334)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient13"
       id="radialGradient14-2"
       cx="43.384182"
       cy="44.199886"
       fx="43.384182"
       fy="44.199886"
       r="41.30278"
       gradientUnits="userSpaceOnUse"
       gradientTransform="translate(60.912832,222.5241)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient1"
       id="radialGradient2-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="translate(53.488946,220.04947)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,95.131459,264.25491)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-94"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,97.300009,287.79051)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-0-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,93.566155,293.51826)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,92.637987,272.87445)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-3-2"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,92.505473,272.13937)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,88.748329,264.91447)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5-88"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,267.44561,122.62379)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,270.7086,127.35093)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-5-5-6"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-46.842714,293.62275)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-8-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,104.92038,270.59533)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-2-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,101.05938,263.23213)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,97.352529,270.98395)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-1-3-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,110.53615,265.73225)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,97.175449,259.20944)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-9-9-6-8-0"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,107.65071,272.14282)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,116.02089,279.52172)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-9-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-170.99192,-240.07837)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-04-5"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,286.80573,-126.51598)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-1-6-9"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-167.73105,-246.71165)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-9-4"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,278.9887,-137.96968)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-2-9-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-267.7689,153.474)" />
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-288.97994,139.58023)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath131">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -253.853,129.20006 -64.67355,-5.42974 26.92803,63.25603 z"
         id="path131" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath141">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -253.853,129.20006 -64.67355,-5.42974 26.92803,63.25603 z"
         id="path141" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath148">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m 264.99289,-104.4642 63.86367,11.557732 -20.78814,-65.530892 z"
         id="path148" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath151">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -152.44278,-240.61421 -0.66083,-64.89772 -60.45116,32.74296 z"
         id="path151" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath154">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m 264.99289,-104.4642 63.86367,11.557732 -20.78814,-65.530892 z"
         id="path154" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath162">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -152.44278,-240.61421 -0.66083,-64.89772 -60.45116,32.74296 z"
         id="path162" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath166">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path166" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath170">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path170" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath174">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path174" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath175">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path175" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath177">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path177" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath178">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path178" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath180">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path180" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath182">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -33.813662,282.82616 -40.482399,50.72795 67.5465585,12.80264 z"
         id="path182" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath183">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m 264.03994,106.84994 38.32633,52.37597 30.08,-61.819404 z"
         id="path183" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath184">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m 264.03994,106.84994 38.32633,52.37597 30.08,-61.819404 z"
         id="path184" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath187">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path187" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath189">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path189" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath190">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path190" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath194">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path194" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath201">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path201" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath210">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path210" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath212">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path212" />
    </clipPath>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath213">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path213" />
    </clipPath>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient214"
       id="radialGradient2-7-2-0-3-7-9-3"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,111.80884,284.75366)" />
    <linearGradient
       id="linearGradient214"
       inkscape:collect="always">
      <stop
         style="stop-color:#b10220;stop-opacity:0.58146107;"
         offset="0"
         id="stop213" />
      <stop
         style="stop-color:#590014;stop-opacity:0.80780524;"
         offset="1"
         id="stop214" />
    </linearGradient>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath198-0">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path198-4" />
    </clipPath>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-4-0-1"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,108.3805,289.60187)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath199-8">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path199-3" />
    </clipPath>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-285.12117,141.68575)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath132-4">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -253.853,129.20006 -64.67355,-5.42974 26.92803,63.25603 z"
         id="path132-1" />
    </clipPath>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient4"
       id="radialGradient2-7-2-2-93-4-87-0-83"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="matrix(0.0710294,0,0,0.0710294,-41.024815,297.58692)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath181-8">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m -33.813662,282.82616 -40.482399,50.72795 67.5465585,12.80264 z"
         id="path181-4" />
    </clipPath>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-8"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-0" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-5"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-1" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-1"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-17" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-16"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-6" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-0"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-8" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-7"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-5" />
    </marker>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-0-6"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-8-0" />
    </marker>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient1"
       id="radialGradient2-8-8"
       cx="50.836403"
       cy="46.676163"
       fx="50.836403"
       fy="46.676163"
       r="37.446667"
       gradientUnits="userSpaceOnUse"
       gradientTransform="translate(53.488946,220.04947)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath212-2">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path212-4" />
    </clipPath>
    <radialGradient
       inkscape:collect="always"
       xlink:href="#linearGradient13"
       id="radialGradient14-2-7"
       cx="43.384182"
       cy="44.199886"
       fx="43.384182"
       fy="44.199886"
       r="41.30278"
       gradientUnits="userSpaceOnUse"
       gradientTransform="translate(60.912832,222.5241)" />
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath213-71">
      <path
         style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:none;stroke-width:1.25979;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="M 104.64827,264.92025 93.134912,328.79194 158.65135,307.95828 Z"
         id="path213-3" />
    </clipPath>
    <marker
       style="overflow:visible"
       id="ConcaveTriangle-9-0-6-8"
       refX="0"
       refY="0"
       orient="auto-start-reverse"
       inkscape:stockid="Concave triangle arrow"
       markerWidth="0.60000002"
       markerHeight="0.60000002"
       viewBox="0 0 1 1"
       inkscape:isstock="true"
       inkscape:collect="always"
       preserveAspectRatio="xMidYMid">
      <path
         transform="scale(0.7)"
         d="M -2,-4 9,0 -2,4 c 2,-2.33 2,-5.66 0,-8 z"
         style="fill:context-stroke;fill-rule:evenodd;stroke:none"
         id="path7-7-8-0-7" />
    </marker>
    <clipPath
       clipPathUnits="userSpaceOnUse"
       id="clipPath237">
      <path
         style="opacity:1;fill:none;fill-opacity:0.972549;fill-rule:evenodd;stroke:#000000;stroke-width:0.750001;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.50001, 4.50001;stroke-dashoffset:0;stroke-opacity:0.960784;paint-order:fill markers stroke"
         d="m 44.012831,95.896295 c 0,0 -6.829845,8.207245 -11.212425,11.125045 -2.439319,1.62402 -8.120293,3.36904 -8.120293,3.36904 l 12.755772,51.97475 37.026653,-42.57425 z"
         id="path237"
         sodipodi:nodetypes="cacccc" />
    </clipPath>
  </defs>
  <g
     inkscape:label="Layer 1"
     inkscape:groupmode="layer"
     id="layer1"
     transform="translate(12.2298,11.2953)">
    <circle
       style="display:inline;fill:#ffffff;fill-opacity:0.803922;fill-rule:evenodd;stroke:url(#radialGradient14);stroke-width:3.9726;stroke-linecap:round;stroke-linejoin:round;paint-order:fill markers stroke"
       id="path9"
       cx="43.384182"
       cy="44.199886"
       r="39.316479" />
    <circle
       style="fill:url(#radialGradient2);fill-rule:evenodd;stroke:none;stroke-width:5.51607;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1"
       cx="43.412518"
       cy="44.201534"
       r="37.446667" />
    <circle
       style="fill:url(#radialGradient2-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2"
       cx="31.092604"
       cy="38.895687"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6"
       cx="37.829502"
       cy="45.046185"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92"
       cx="34.194386"
       cy="38.011673"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92-1"
       cx="45.246918"
       cy="73.908669"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62-0-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92-1-9"
       cx="35.979851"
       cy="13.810245"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62-0-9-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92-1-9-0"
       cx="70.79023"
       cy="49.037834"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62-0-9-5-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92-1-9-0-5"
       cx="14.005543"
       cy="38.352364"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-62-0-9-5-9-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-92-1-9-0-5-9"
       cx="63.513981"
       cy="49.491066"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44"
       cx="23.853704"
       cy="40.593117"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6"
       cx="25.17919"
       cy="62.865765"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1"
       cx="39.998074"
       cy="68.581779"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-4-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-6-5"
       cx="51.078564"
       cy="70.393143"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8"
       cx="53.977749"
       cy="66.603271"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3"
       cx="26.454466"
       cy="33.242321"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8"
       cx="61.781498"
       cy="47.054893"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3"
       cx="27.960974"
       cy="69.937691"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-0"
       cx="36.264229"
       cy="74.30954"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9"
       cx="19.739368"
       cy="52.140484"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9"
       cx="26.649704"
       cy="56.592941"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9-8"
       cx="42.235508"
       cy="70.911507"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9-8-8"
       cx="35.336079"
       cy="53.665718"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9-8-8-4"
       cx="35.203564"
       cy="52.930649"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-4"
       cx="34.353489"
       cy="32.262413"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9"
       cx="31.446379"
       cy="45.70575"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5"
       cx="26.630733"
       cy="53.269852"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8"
       cx="18.042452"
       cy="60.42112"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2"
       cx="67.878929"
       cy="16.640438"
       r="2.6598144"
       transform="rotate(46.413219)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2"
       cx="71.14193"
       cy="21.36758"
       r="2.6598144"
       transform="rotate(46.413219)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2-9"
       cx="8.9167852"
       cy="72.198555"
       r="2.6598144"
       transform="rotate(-28.372626)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2-1"
       cx="11.791796"
       cy="79.384583"
       r="2.6598144"
       transform="rotate(-28.372626)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-9"
       cx="47.618443"
       cy="50.857445"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-8-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-9-6"
       cx="46.409824"
       cy="39.041035"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-2"
       cx="43.757427"
       cy="44.023403"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29"
       cx="40.050579"
       cy="51.775234"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-7"
       cx="52.554768"
       cy="55.326233"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-1-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-7-9"
       cx="53.234211"
       cy="46.523525"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5"
       cx="39.873493"
       cy="40.000717"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-8"
       cx="54.785801"
       cy="38.476456"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-0"
       cx="44.252659"
       cy="31.559181"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-2"
       cx="13.797639"
       cy="41.837181"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-6-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-2-7"
       cx="49.290405"
       cy="57.167439"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-6-8-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-2-7-2"
       cx="23.691412"
       cy="65.034996"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7"
       cx="21.30097"
       cy="48.690395"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3"
       cx="57.131485"
       cy="60.842175"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1"
       cx="-20.690973"
       cy="54.218403"
       r="2.6598144"
       transform="rotate(-82.959297)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1-6"
       cx="16.824659"
       cy="43.77985"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1-6-7"
       cx="20.240057"
       cy="35.625771"
       r="2.6598144" />
    <circle
       style="fill:url(#radialGradient2-7-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-9"
       cx="-65.844269"
       cy="-29.597292"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-1"
       cx="-59.107365"
       cy="-23.446787"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-38);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-0"
       cx="-73.083168"
       cy="-27.899858"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-7"
       cx="54.413609"
       cy="-16.220074"
       r="2.6598144"
       transform="rotate(89.960195)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-5"
       cx="-44.133724"
       cy="-12.767736"
       r="2.6598144"
       transform="rotate(-167.54011)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-8"
       cx="30.710732"
       cy="30.892342"
       r="2.6598144"
       transform="rotate(-7.9910847)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-64);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-7"
       cx="-32.515396"
       cy="-41.445763"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-0"
       cx="-32.752232"
       cy="21.438061"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-04);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-4"
       cx="67.848808"
       cy="-60.325703"
       r="2.6598144"
       transform="rotate(89.960195)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-0-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-0-8"
       cx="-47.867573"
       cy="-7.0399833"
       r="2.6598144"
       transform="rotate(-167.54011)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-0"
       cx="24.501656"
       cy="25.067587"
       r="2.6598144"
       transform="rotate(-7.9910847)" />
    <circle
       style="fill:url(#radialGradient2-7-2-1-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-4-4"
       cx="-62.583378"
       cy="-36.23056"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-296"
       cx="-65.490494"
       cy="-22.787226"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-56);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-1"
       cx="-70.306137"
       cy="-15.223124"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-0"
       transform="rotate(89.960195)"
       r="2.6598144"
       cy="-73.030563"
       cx="62.048859" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2-4"
       cx="-48.566013"
       cy="39.632168"
       r="2.6598144"
       transform="rotate(-122.78511)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2-2"
       cx="-45.786922"
       cy="26.220222"
       r="2.6598144"
       transform="rotate(-121.12689)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5-5-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2-9-2"
       cx="23.56934"
       cy="-42.515446"
       r="2.6598144"
       transform="rotate(79.469743)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87-0-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2-1-2"
       cx="11.835324"
       cy="36.644485"
       r="2.6598144"
       transform="rotate(-36.363714)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-8-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-9-0"
       cx="26.448578"
       cy="19.684523"
       r="2.6598144"
       transform="rotate(-7.9910847)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-8-6-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-9-6-5"
       cx="-39.158039"
       cy="-0.34544733"
       r="2.6598144"
       transform="rotate(-128.44305)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-2"
       cx="-1.5695429"
       cy="-56.121792"
       r="2.6598144"
       transform="rotate(107.84237)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-1-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-7-90"
       cx="32.435329"
       cy="21.908049"
       r="2.6598144"
       transform="rotate(-7.9910847)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-1-3-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-7-9-2"
       cx="24.22644"
       cy="31.13665"
       r="2.6598144"
       transform="rotate(-7.9910847)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-7);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-83"
       cx="-57.063374"
       cy="-28.492258"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-5-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-8-8"
       cx="-30.782063"
       cy="-0.91003013"
       r="2.6598144"
       transform="rotate(-128.44305)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-1-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-0-0"
       cx="-49.498684"
       cy="68.154778"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-6-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-2-4"
       cx="-64.239456"
       cy="-16.250299"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-0"
       cx="-75.635902"
       cy="-19.802576"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9"
       cx="-65.733444"
       cy="63.344986"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9-1"
       cx="-69.592209"
       cy="61.239464"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9-1-4"
       cx="-18.609303"
       cy="67.750542"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-0-4);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9-1-4-8"
       cx="-50.284912"
       cy="18.309175"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1-1"
       cx="-18.602438"
       cy="55.612053"
       r="2.6598144"
       transform="rotate(-84.580811)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-8-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1-6-7-6"
       cx="-76.696815"
       cy="-32.867195"
       r="2.6598144"
       transform="rotate(-169.19833)" />
    <g
       id="g19"
       transform="translate(22.378079,47.944485)">
      <rect
         style="fill:#ffffff;fill-rule:evenodd;stroke:none;stroke-width:0.3;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         id="rect24"
         width="1.8138908"
         height="2.4575295"
         x="70.085442"
         y="80.768097"
         transform="rotate(-54.146651)" />
      <g
         id="g21"
         transform="matrix(1.4367106,0,0,1.4367106,-72.171108,-2.2943584)">
        <circle
           style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-4);fill-rule:evenodd;stroke:none;stroke-width:1.53352;stroke-linecap:round;paint-order:fill markers stroke"
           id="path1-2-6-44-6-1-8-3-8-3-7-3-7"
           cx="126.30329"
           cy="-11.762299"
           r="10.410519" />
        <path
           style="fill:#a05a2c;fill-rule:evenodd;stroke:#a05a2c;stroke-width:0.439317;stroke-linecap:round;stroke-dasharray:2.6359, 2.6359;stroke-dashoffset:0;paint-order:fill markers stroke"
           d="M 138.10398,-26.510674 V -3.8151456"
           id="path8" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:#4d4d4d;stroke-width:0.443095;stroke-linecap:round;stroke-dasharray:0.886192, 0.886192;stroke-dashoffset:0;marker-start:url(#ArrowWide);paint-order:fill markers stroke"
           d="m 125.92215,-28.515815 v 16.96846"
           id="path8-9" />
        <path
           style="fill:#a05a2c;fill-rule:evenodd;stroke:#a05a2c;stroke-width:0.476627;stroke-linecap:round;stroke-dasharray:2.85974, 2.85974;stroke-dashoffset:0;paint-order:fill markers stroke"
           d="m 125.88481,-11.571508 13.18796,8.3783534"
           id="path8-6" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:#4d4d4d;stroke-width:0.425331;stroke-linecap:round;stroke-dasharray:0.850662, 0.850662;stroke-dashoffset:0;marker-end:url(#marker14-7);paint-order:fill markers stroke"
           d="m 125.9152,-11.600949 19.19958,4.5829924"
           id="path8-6-8" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:#4d4d4d;stroke-width:0.525022;stroke-linecap:round;stroke-dasharray:1.05005, 1.05005;stroke-dashoffset:0;marker-end:url(#marker13);paint-order:fill markers stroke"
           d="M 125.82182,-11.48688 113.4786,-2.9294186"
           id="path8-6-9" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:url(#linearGradient7);stroke-width:0.926954;stroke-linecap:round;stroke-dasharray:none;marker-end:url(#ConcaveTriangle);paint-order:fill markers stroke"
           d="m 126.24026,-11.820421 9.73244,-12.069217"
           id="path4"
           sodipodi:nodetypes="cc" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:#552200;stroke-width:0.395302;stroke-linecap:round;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
           id="path11-6"
           sodipodi:type="arc"
           sodipodi:cx="31.582554"
           sodipodi:cy="-134.427"
           sodipodi:rx="16.341784"
           sodipodi:ry="13.513863"
           sodipodi:start="0"
           sodipodi:end="0.69025833"
           sodipodi:open="true"
           sodipodi:arc-type="arc"
           d="m 47.924337,-134.427 a 16.341784,13.513863 0 0 1 -3.740935,8.60477"
           transform="matrix(0.16581651,0.98615662,-0.91086531,0.41270375,0,0)" />
        <path
           style="fill:none;fill-rule:evenodd;stroke:#552200;stroke-width:0.406833;stroke-linecap:round;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
           id="path11-6-6"
           sodipodi:type="arc"
           sodipodi:cx="-0.63133687"
           sodipodi:cy="125.6298"
           sodipodi:rx="8.4097376"
           sodipodi:ry="6.9544449"
           sodipodi:start="0"
           sodipodi:end="0.69025833"
           sodipodi:open="true"
           sodipodi:arc-type="arc"
           d="m 7.7784007,125.6298 a 8.4097376,6.9544449 0 0 1 -1.9251441,4.42815"
           transform="matrix(0.16236497,-0.98673077,0.99541971,-0.09560129,0,0)" />
        <g
           transform="matrix(0.40183383,0,0,0.40183383,126.73953,-18.369524)"
           ns58:version="1.11.1"
           ns58:texconverter="pdflatex"
           ns58:pdfconverter="inkscape"
           ns58:text="$\\theta$"
           ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
           ns58:scale="2.441120244458815"
           ns58:alignment="middle center"
           ns58:inkscapeversion="1.4.2"
           ns58:jacobian_sqrt="0.861174"
           id="g15"
           style="fill:#502d16;stroke-width:2;stroke-dasharray:none">
          <defs
             id="id-dfeafae5-ced4-450b-99dd-714855df862c" />
          <g
             fill="#000000"
             fill-opacity="1"
             id="id-2419b262-1e83-4f7e-aca8-4eb59131b1a6"
             transform="translate(-149.134,-127.734)"
             style="fill:#502d16;stroke-width:2;stroke-dasharray:none">
            <g
               transform="translate(148.712,134.765)"
               id="g14"
               style="fill:#502d16;stroke-width:2;stroke-dasharray:none">
              <path
                 d="m 4.53125,-4.984375 c 0,-0.65625 -0.171875,-2.046875 -1.1875,-2.046875 -1.390625,0 -2.921875,2.8125 -2.921875,5.09375 0,0.9375 0.28125,2.046875 1.1875,2.046875 1.40625,0 2.921875,-2.859375 2.921875,-5.09375 z M 1.46875,-3.625 C 1.640625,-4.25 1.84375,-5.046875 2.25,-5.765625 2.515625,-6.25 2.875,-6.8125 3.328125,-6.8125 c 0.484375,0 0.546875,0.640625 0.546875,1.203125 0,0.5 -0.078125,1 -0.3125,1.984375 z m 2,0.328125 C 3.359375,-2.84375 3.15625,-2 2.765625,-1.28125 c -0.34375,0.6875 -0.71875,1.171875 -1.15625,1.171875 -0.328125,0 -0.53125,-0.296875 -0.53125,-1.21875 0,-0.421875 0.0625,-1 0.3125,-1.96875 z m 0,0"
                 id="id-7dace4ee-b2dc-4a8d-ad48-35f4897792fa"
                 style="fill:#502d16;stroke-width:2;stroke-dasharray:none" />
            </g>
          </g>
        </g>
        <g
           transform="matrix(0.40183365,0,0,0.40183365,124.78358,-5.8026556)"
           ns58:version="1.11.1"
           ns58:texconverter="pdflatex"
           ns58:pdfconverter="inkscape"
           ns58:text="$\\varphi$"
           ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
           ns58:scale="1.3008661053983923"
           ns58:alignment="middle center"
           ns58:inkscapeversion="1.4.2"
           ns58:jacobian_sqrt="0.458917"
           style="fill:#502d16;stroke:#502d16;stroke-width:0"
           id="g18">
          <defs
             id="id-a44466a7-9a38-47c6-b9b7-23e2b48a4409"
             style="fill:#502d16;stroke-width:0" />
          <g
             fill-opacity="1"
             id="id-0e1852ba-b304-414f-b6ae-83f3b4ffac72"
             transform="translate(-149.212,-130.359)"
             style="fill:#502d16;stroke:#502d16;stroke-width:0">
            <g
               transform="translate(148.712,134.765)"
               style="fill:#502d16;stroke:#502d16;stroke-width:0"
               id="g17">
              <path
                 d="M 1.6875,1.6875 C 1.65625,1.828125 1.640625,1.84375 1.640625,1.890625 c 0,0.21875 0.1875,0.28125 0.296875,0.28125 0.046875,0 0.265625,-0.03125 0.359375,-0.265625 C 2.328125,1.828125 2.375,1.5 2.65625,0.09375 c 0.078125,0 0.15625,0.015625 0.328125,0.015625 1.65625,0 3.1875,-1.5625 3.1875,-3.140625 0,-0.78125 -0.390625,-1.375 -1.140625,-1.375 -1.4375,0 -2.046875,1.9375 -2.640625,3.875 C 1.3125,-0.734375 0.75,-1.28125 0.75,-2 c 0,-0.28125 0.234375,-1.375 0.828125,-2.0625 0.09375,-0.09375 0.09375,-0.109375 0.09375,-0.140625 0,-0.03125 -0.03125,-0.09375 -0.125,-0.09375 -0.28125,0 -1.046875,1.453125 -1.046875,2.40625 0,0.9375 0.65625,1.65625 1.71875,1.90625 z m 1.390625,-2.15625 c -0.09375,0 -0.109375,0 -0.1875,-0.015625 -0.125,0 -0.125,0 -0.125,-0.03125 0,-0.015625 0.171875,-0.9375 0.1875,-1.078125 0.3125,-1.28125 1.09375,-2.234375 1.984375,-2.234375 0.6875,0 0.953125,0.53125 0.953125,1.015625 0,1.125 -1.28125,2.34375 -2.8125,2.34375 z m 0,0"
                 id="id-901225e4-231d-4c15-9a15-8cef40283c59"
                 style="fill:#502d16;stroke:#502d16;stroke-width:0" />
            </g>
          </g>
        </g>
      </g>
      <text
         xml:space="preserve"
         style="font-size:3.175px;font-family:'DejaVu Sans';-inkscape-font-specification:'DejaVu Sans';text-align:center;writing-mode:lr-tb;direction:ltr;text-anchor:middle;fill:#a05a2c;fill-rule:evenodd;stroke:#a05a2c;stroke-width:0.4;stroke-linecap:round;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         x="96.180817"
         y="-12.21375"
         id="text19"><tspan
           sodipodi:role="line"
           id="tspan19"
           style="stroke-width:0.4"
           x="96.180817"
           y="-12.21375" /></text>
      <g
         transform="matrix(0.57943596,0,0,0.57943596,115.69858,-44.902021)"
         ns58:version="1.11.1"
         ns58:texconverter="pdflatex"
         ns58:pdfconverter="inkscape"
         ns58:text="$\\mathbf{F_a}$"
         ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
         ns58:scale="1.3008661053983923"
         ns58:alignment="middle center"
         ns58:inkscapeversion="1.4.2"
         ns58:jacobian_sqrt="0.458917"
         id="g24">
        <defs
           id="id-0bbeb6e6-5e62-4704-8bdc-f568b397a3f8" />
        <g
           fill="#000000"
           fill-opacity="1"
           id="id-33328e6d-c650-42d1-8402-3102d0ec786c"
           transform="translate(-149.103,-127.984)">
          <g
             transform="translate(148.712,134.765)"
             id="g22">
            <path
               d="M 6.421875,-6.78125 H 0.390625 V -6.3125 H 1.46875 v 5.84375 H 0.390625 V 0 c 0.375,-0.03125 1.390625,-0.03125 1.828125,-0.03125 0.484375,0 1.5625,0 2.015625,0.03125 V -0.46875 H 2.875 v -2.6875 h 0.5 c 0.96875,0 1.046875,0.421875 1.046875,1.15625 h 0.46875 V -4.796875 H 4.421875 C 4.421875,-4.0625 4.34375,-3.625 3.375,-3.625 h -0.5 v -2.6875 h 1.40625 c 1.59375,0 1.828125,0.765625 1.984375,1.9375 h 0.46875 z m 0,0"
               id="id-2e43cc0c-40ae-461d-b2f0-a03cc3a495c0" />
          </g>
        </g>
        <g
           fill="#000000"
           fill-opacity="1"
           id="id-a2559208-40c1-4e50-ad16-18953353bfed"
           transform="translate(-149.103,-127.984)">
          <g
             transform="translate(155.921,136.259)"
             id="g23">
            <path
               d="m 3.671875,-2.0625 c 0,-0.5625 -0.453125,-1.09375 -1.703125,-1.09375 -0.40625,0 -1.390625,0 -1.390625,0.6875 0,0.3125 0.234375,0.484375 0.484375,0.484375 0.3125,0 0.484375,-0.203125 0.484375,-0.46875 0,-0.15625 -0.0625,-0.265625 -0.078125,-0.28125 -0.015625,-0.03125 -0.015625,-0.046875 -0.015625,-0.046875 0,-0.046875 0.4375,-0.0625 0.484375,-0.0625 0.5,0 0.859375,0.203125 0.859375,0.796875 v 0.1875 c -0.34375,0 -2.515625,0.03125 -2.515625,1.0625 0,0.640625 0.765625,0.84375 1.46875,0.84375 0.734375,0 1.0625,-0.34375 1.1875,-0.515625 C 2.9375,-0.171875 3.125,0 3.6875,0 h 0.421875 c 0.125,0 0.234375,0 0.234375,-0.1875 0,-0.203125 -0.09375,-0.203125 -0.25,-0.203125 -0.421875,0 -0.421875,-0.0625 -0.421875,-0.21875 z m -0.875,1.109375 c 0,0.140625 0,0.34375 -0.28125,0.515625 -0.25,0.15625 -0.578125,0.15625 -0.625,0.15625 C 1.5,-0.28125 1.15625,-0.5 1.15625,-0.8125 c 0,-0.5625 0.9375,-0.75 1.640625,-0.78125 z m 0,0"
               id="id-116be6f9-33a3-4d03-9a69-c4029460aaec" />
          </g>
        </g>
      </g>
      <g
         transform="matrix(0.57645496,-0.05870061,0.05870061,0.57645496,102.75354,28.653901)"
         ns58:version="1.11.1"
         ns58:texconverter="pdflatex"
         ns58:pdfconverter="inkscape"
         ns58:text="$\\mathbf{F_m}$"
         ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
         ns58:scale="1.6424943957468967"
         ns58:alignment="middle center"
         ns58:inkscapeversion="1.4.2"
         ns58:jacobian_sqrt="0.579436"
         id="g24-2"
         style="fill:#ffffff">
        <defs
           id="id-64b6a99a-3003-4bb6-8fcc-28ec40724c25" />
        <g
           fill="#000000"
           fill-opacity="1"
           id="id-3205149d-ceb4-4529-9829-afb16aa74cf2"
           transform="translate(-149.103,-127.984)"
           style="fill:#ffffff">
          <g
             transform="translate(148.712,134.765)"
             id="g32"
             style="fill:#ffffff">
            <path
               d="M 6.421875,-6.78125 H 0.390625 V -6.3125 H 1.46875 v 5.84375 H 0.390625 V 0 c 0.375,-0.03125 1.390625,-0.03125 1.828125,-0.03125 0.484375,0 1.5625,0 2.015625,0.03125 V -0.46875 H 2.875 v -2.6875 h 0.5 c 0.96875,0 1.046875,0.421875 1.046875,1.15625 h 0.46875 V -4.796875 H 4.421875 C 4.421875,-4.0625 4.34375,-3.625 3.375,-3.625 h -0.5 v -2.6875 h 1.40625 c 1.59375,0 1.828125,0.765625 1.984375,1.9375 h 0.46875 z m 0,0"
               id="id-f3275edb-d225-46f2-9500-3e39318f18ab"
               style="fill:#ffffff" />
          </g>
        </g>
        <g
           fill="#000000"
           fill-opacity="1"
           id="id-e3c8fcf3-ea61-4d4d-bf30-5f029a7e587d"
           transform="translate(-149.103,-127.984)"
           style="fill:#ffffff">
          <g
             transform="translate(155.921,136.259)"
             id="g33"
             style="fill:#ffffff">
            <path
               d="m 6.75,-2.09375 c 0,-0.875 -0.578125,-1.046875 -1.203125,-1.046875 -0.65625,0 -1.09375,0.3125 -1.3125,0.65625 -0.171875,-0.609375 -0.78125,-0.65625 -1.15625,-0.65625 -0.828125,0 -1.234375,0.5 -1.375,0.734375 v -0.734375 l -1.25,0.0625 V -2.6875 c 0.40625,0 0.453125,0 0.453125,0.265625 v 2.03125 H 0.453125 V 0 c 0,0 0.5625,-0.03125 0.90625,-0.03125 C 1.6875,-0.03125 2.265625,0 2.265625,0 v -0.390625 h -0.46875 v -1.34375 c 0,-0.828125 0.75,-1.078125 1.140625,-1.078125 0.3125,0 0.453125,0.15625 0.453125,0.671875 v 1.75 H 2.921875 V 0 c 0,0 0.5625,-0.03125 0.90625,-0.03125 0.34375,0 0.90625,0.03125 0.90625,0.03125 v -0.390625 h -0.46875 v -1.34375 c 0,-0.828125 0.75,-1.078125 1.15625,-1.078125 0.3125,0 0.4375,0.15625 0.4375,0.671875 v 1.75 H 5.390625 V 0 C 5.40625,0 5.96875,-0.03125 6.296875,-0.03125 6.640625,-0.03125 7.203125,0 7.21875,0 V -0.390625 H 6.75 Z m 0,0"
               id="id-afd02088-cb65-432f-aa92-096a7618dd19"
               style="fill:#ffffff" />
          </g>
        </g>
      </g>
      <path
         style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         d="M 53.003783,-12.61078 101.49315,-33.702353"
         id="path21"
         sodipodi:nodetypes="cc" />
      <path
         style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         d="m 53.607339,-5.0244265 51.481771,2.1407144"
         id="path21-0"
         sodipodi:nodetypes="cc" />
      <path
         d="M 66.792353,-5.5956563"
         style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         id="path1-1" />
      <path
         d="M 49.424638,17.391095 89.463841,47.471102"
         style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         id="path1-26"
         sodipodi:nodetypes="cc" />
      <path
         d="M 52.040387,10.796392 98.704382,24.458466"
         style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
         id="path1-4"
         sodipodi:nodetypes="cc" />
    </g>
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-0-8-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-1-6-9"
       cx="-80.112213"
       cy="-24.713129"
       r="2.6598144"
       transform="rotate(-169.19833)"
       inkscape:label="path1-2-6-44-6-1-8-3-8-3-7-3-1-6-9" />
    <circle
       style="display:inline;fill:#ffffff;fill-opacity:0.803922;fill-rule:evenodd;stroke:url(#radialGradient14-2);stroke-width:3.9726;stroke-linecap:round;stroke-linejoin:round;paint-order:fill markers stroke"
       id="path9-4"
       cx="104.29701"
       cy="266.724"
       r="39.316479"
       clip-path="url(#clipPath213)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-8);fill-rule:evenodd;stroke:none;stroke-width:5.51607;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-9"
       cx="104.32535"
       cy="266.72565"
       r="37.446667"
       clip-path="url(#clipPath212)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <g
       id="g233"
       transform="matrix(0.94943619,-0.67245706,0.67245706,0.94943619,11.074771,2.1603721)"
       clip-path="url(#clipPath237)">
      <circle
         style="display:inline;fill:#ffffff;fill-opacity:0.803922;fill-rule:evenodd;stroke:url(#radialGradient14-2-7);stroke-width:3.9726;stroke-linecap:round;stroke-linejoin:round;paint-order:fill markers stroke"
         id="path9-4-8"
         cx="104.29701"
         cy="266.724"
         r="39.316479"
         clip-path="url(#clipPath213-71)"
         transform="matrix(1.3133802,0,0,1.3133802,-118.44171,-261.00389)" />
      <circle
         style="fill:url(#radialGradient2-8-8);fill-rule:evenodd;stroke:none;stroke-width:5.51607;stroke-linecap:round;paint-order:fill markers stroke"
         id="path1-9-5"
         cx="104.32535"
         cy="266.72565"
         r="37.446667"
         clip-path="url(#clipPath212-2)"
         transform="matrix(1.3133802,0,0,1.3133802,-118.44171,-261.00389)" />
    </g>
    <circle
       style="fill:url(#radialGradient2-7-2-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-5"
       cx="98.742332"
       cy="267.57028"
       r="2.6598144"
       clip-path="url(#clipPath210)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-94);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-57"
       cx="100.9109"
       cy="291.10587"
       r="2.6598144"
       clip-path="url(#clipPath201)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-0-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-0-2"
       cx="97.177063"
       cy="296.83365"
       r="2.6598144"
       clip-path="url(#clipPath194)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9-8-8-9"
       cx="96.248909"
       cy="276.18982"
       r="2.6598144"
       clip-path="url(#clipPath190)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-2-4-2-2-3-2);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-9-9-8-8-4-0"
       cx="96.116394"
       cy="275.45474"
       r="2.6598144"
       clip-path="url(#clipPath189)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-0"
       cx="92.359215"
       cy="268.22986"
       r="2.6598144"
       clip-path="url(#clipPath187)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5-88);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2-2"
       cx="271.05652"
       cy="125.93917"
       r="2.6598144"
       transform="matrix(0.90551318,0.95132191,-0.95132191,0.90551318,-68.92316,-244.01494)"
       clip-path="url(#clipPath184)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2-12"
       cx="274.31952"
       cy="130.66632"
       r="2.6598144"
       transform="matrix(0.90551318,0.95132191,-0.95132191,0.90551318,-68.92316,-244.01494)"
       clip-path="url(#clipPath183)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-5-5-6);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-2-9-0"
       cx="-43.231812"
       cy="296.93811"
       r="2.6598144"
       transform="matrix(1.1556113,-0.62412337,0.62412337,1.1556113,-68.923156,-244.01494)"
       clip-path="url(#clipPath182)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-8-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-9-3"
       cx="108.53127"
       cy="273.91071"
       r="2.6598144"
       clip-path="url(#clipPath180)"
       transform="matrix(1.3133802,0,0,1.3133802,-71.342798,-242.74749)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-2-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-2-1"
       cx="104.67026"
       cy="266.54752"
       r="2.6598144"
       clip-path="url(#clipPath178)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-9"
       cx="100.96341"
       cy="274.29935"
       r="2.6598144"
       clip-path="url(#clipPath177)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-1-3-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-7-9-5"
       cx="114.14704"
       cy="269.04764"
       r="2.6598144"
       clip-path="url(#clipPath175)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-4);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-6"
       cx="100.78632"
       cy="262.52481"
       r="2.6598144"
       clip-path="url(#clipPath174)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-9-9-6-8-0);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-29-5-2-7-6"
       cx="111.26157"
       cy="275.45819"
       r="2.6598144"
       clip-path="url(#clipPath170)"
       transform="matrix(1.3133802,0,0,1.3133802,-70.510657,-247.18994)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-8"
       cx="119.63183"
       cy="282.8371"
       r="2.6598144"
       clip-path="url(#clipPath166)"
       transform="matrix(1.3133802,0,0,1.3133802,-68.923156,-244.01492)" />
    <circle
       style="fill:url(#radialGradient2-7-9-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-9-6"
       cx="-167.38106"
       cy="-236.76299"
       r="2.6598144"
       transform="matrix(-1.2901094,-0.24614051,0.24614051,-1.2901094,-68.923156,-244.01493)"
       clip-path="url(#clipPath162)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-04-5);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-4-9"
       cx="290.41663"
       cy="-123.2006"
       r="2.6598144"
       transform="matrix(9.1244231e-4,1.3133799,-1.3133799,9.1244231e-4,-68.923156,-244.01493)"
       clip-path="url(#clipPath154)" />
    <circle
       style="fill:url(#radialGradient2-7-2-1-6-9);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-4-4-7"
       cx="-164.12018"
       cy="-243.39626"
       r="2.6598144"
       transform="matrix(-1.2901094,-0.24614051,0.24614051,-1.2901094,-68.923156,-244.01493)"
       clip-path="url(#clipPath151)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-9-4);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-0-0"
       transform="matrix(9.1244231e-4,1.3133799,-1.3133799,9.1244231e-4,-71.777993,-249.98413)"
       r="2.6598144"
       cy="-134.6543"
       cx="282.59958"
       clip-path="url(#clipPath148)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-2-9-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-2-5-4"
       cx="-264.15802"
       cy="156.78938"
       r="2.6598144"
       transform="matrix(0.1240379,-1.3075099,1.3075099,0.1240379,-68.923156,-244.01494)"
       clip-path="url(#clipPath141)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-1-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9-1-5"
       cx="-285.36899"
       cy="142.8956"
       r="2.6598144"
       transform="matrix(0.1240379,-1.3075099,1.3075099,0.1240379,-68.923156,-244.01494)"
       clip-path="url(#clipPath131)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-9-7);fill-rule:evenodd;stroke:none;stroke-width:1.01801;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-0-9"
       transform="rotate(105.4693)"
       r="6.9108567"
       cy="-155.39909"
       cx="50.918571" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-8);paint-order:fill markers stroke"
       d="m 88.309634,127.31553 2.225888,1.74518"
       id="path35-7-9"
       sodipodi:nodetypes="cc" />
    <g
       transform="matrix(0.75868569,0.00674141,-0.00674141,0.75868569,145.43188,94.837952)"
       ns58:version="1.11.1"
       ns58:texconverter="pdflatex"
       ns58:pdfconverter="inkscape"
       ns58:text="$\\nabla\\phi$"
       ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
       ns58:scale="1.6424943957468967"
       ns58:alignment="middle center"
       ns58:inkscapeversion="1.4.2"
       ns58:jacobian_sqrt="0.579436"
       id="g38"
       style="fill:#800000;stroke:none">
      <defs
         id="id-aa40f5b1-5a85-4c3a-af8f-9fed8d09de9f" />
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-90caa7c7-814f-40f8-93b7-dd90eea1d04a"
         transform="translate(-149.181,-127.843)"
         style="fill:#800000;stroke:none">
        <g
           transform="translate(148.712,134.765)"
           id="g36"
           style="fill:#800000;stroke:none">
          <path
             d="M 7.78125,-6.59375 C 7.796875,-6.625 7.828125,-6.6875 7.828125,-6.734375 7.828125,-6.796875 7.8125,-6.8125 7.59375,-6.8125 H 0.703125 c -0.21875,0 -0.234375,0.015625 -0.234375,0.078125 0,0.046875 0.03125,0.109375 0.046875,0.140625 L 3.875,0.140625 c 0.078125,0.125 0.109375,0.1875 0.265625,0.1875 0.171875,0 0.203125,-0.0625 0.28125,-0.1875 z m -6.078125,0.5 h 5.46875 l -2.71875,5.484375 z m 0,0"
             id="id-c1a9057d-1119-4e11-b38e-e9746b08c735"
             style="fill:#800000;stroke:none" />
        </g>
      </g>
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-be637cfa-0d5f-46d3-ba9a-a15d12ec3353"
         transform="translate(-149.181,-127.843)"
         style="fill:#800000;stroke:none">
        <g
           transform="translate(157.014,134.765)"
           id="g37"
           style="fill:#800000;stroke:none">
          <path
             d="m 4.359375,-6.671875 c 0,-0.03125 0.03125,-0.140625 0.03125,-0.140625 0,-0.015625 0,-0.109375 -0.125,-0.109375 -0.09375,0 -0.109375,0.03125 -0.15625,0.203125 L 3.53125,-4.421875 c -1.578125,0.0625 -3.046875,1.375 -3.046875,2.734375 0,0.953125 0.703125,1.734375 1.921875,1.8125 C 2.328125,0.421875 2.25,0.75 2.171875,1.0625 c -0.125,0.46875 -0.21875,0.84375 -0.21875,0.875 0,0.09375 0.078125,0.109375 0.125,0.109375 C 2.125,2.046875 2.140625,2.03125 2.171875,2 2.1875,1.984375 2.25,1.75 2.28125,1.609375 L 2.65625,0.125 c 1.609375,-0.0625 3.0625,-1.40625 3.0625,-2.734375 0,-0.796875 -0.53125,-1.703125 -1.921875,-1.8125 z m -1.90625,6.578125 c -0.59375,-0.03125 -1.3125,-0.390625 -1.3125,-1.375 0,-1.203125 0.859375,-2.59375 2.34375,-2.734375 z m 1.28125,-4.109375 c 0.765625,0.046875 1.328125,0.5 1.328125,1.375 0,1.1875 -0.859375,2.609375 -2.34375,2.734375 z m 0,0"
             id="id-10e59b98-cfdc-4242-b699-e57d347961e3"
             style="fill:#800000;stroke:none" />
        </g>
      </g>
    </g>
    <g
       sodipodi:type="inkscape:box3d"
       id="g219"
       style="opacity:1;fill:none;fill-opacity:0.972549;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0;stroke-opacity:0.960784;paint-order:fill markers stroke"
       inkscape:perspectiveID="#perspective219"
       inkscape:corner0="2.2277825 : -0.10703232 : 0 : 1"
       inkscape:corner7="1.770409 : -0.16432786 : 0.15167482 : 1">
      <path
         sodipodi:type="inkscape:box3dside"
         id="path224"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="11"
         d="m 80.919046,122.58123 13.240776,3.72619 v 15.82119 l -13.240776,-3.72618 z"
         points="94.159822,126.30742 94.159822,142.12861 80.919046,138.40243 80.919046,122.58123 " />
      <path
         sodipodi:type="inkscape:box3dside"
         id="path219"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="6"
         d="m 66.746097,125.54686 v 18.22087 l 14.172949,-5.3653 v -15.8212 z"
         points="66.746097,143.76773 80.919046,138.40243 80.919046,122.58123 66.746097,125.54686 " />
      <path
         sodipodi:type="inkscape:box3dside"
         id="path223"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="13"
         d="m 66.746097,143.76773 15.249069,4.29135 12.164656,-5.93047 -13.240776,-3.72618 z"
         points="81.995166,148.05908 94.159822,142.12861 80.919046,138.40243 66.746097,143.76773 " />
      <path
         sodipodi:type="inkscape:box3dside"
         id="path220"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="5"
         d="m 66.746097,125.54686 15.249069,4.29135 12.164656,-3.53079 -13.240776,-3.72619 z"
         points="81.995166,129.83821 94.159822,126.30742 80.919046,122.58123 66.746097,125.54686 " />
      <path
         sodipodi:type="inkscape:box3dside"
         id="path222"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="14"
         d="m 81.995166,129.83821 v 18.22087 l 12.164656,-5.93047 v -15.82119 z"
         points="81.995166,148.05908 94.159822,142.12861 94.159822,126.30742 81.995166,129.83821 " />
      <path
         sodipodi:type="inkscape:box3dside"
         id="path221"
         style="fill:none;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.75;stroke-linecap:butt;stroke-linejoin:bevel;stroke-dasharray:4.5, 4.5;stroke-dashoffset:0"
         inkscape:box3dsidetype="3"
         d="m 66.746097,125.54686 15.249069,4.29135 v 18.22087 l -15.249069,-4.29135 z"
         points="81.995166,129.83821 81.995166,148.05908 66.746097,143.76773 66.746097,125.54686 " />
    </g>
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-3);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-1"
       cx="115.41975"
       cy="288.06903"
       r="2.6598144"
       clip-path="url(#clipPath198-0)"
       transform="matrix(1.5511867,0,0,1.5511867,-98.269893,-311.09202)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-4-0-1);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-6-5-8"
       cx="111.99139"
       cy="292.91724"
       r="2.6598144"
       clip-path="url(#clipPath199-8)"
       transform="matrix(1.3133802,0,0,1.3133802,-69.820123,-244.53152)" />
    <circle
       style="fill:url(#radialGradient2-7-2-0-3-7-9-8-6-7-9-8-1-8);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-44-6-1-8-3-8-3-7-3-9-4"
       cx="-281.51022"
       cy="145.00111"
       r="2.6598144"
       transform="matrix(0.1240379,-1.3075099,1.3075099,0.1240379,-67.427479,-246.05549)"
       clip-path="url(#clipPath132-4)" />
    <circle
       style="fill:url(#radialGradient2-7-2-2-93-4-87-0-83);fill-rule:evenodd;stroke:none;stroke-width:0.391804;stroke-linecap:round;paint-order:fill markers stroke"
       id="path1-2-6-9-5-8-2-1-7"
       cx="-37.413902"
       cy="300.90228"
       r="2.6598144"
       transform="matrix(1.1556113,-0.62412337,0.62412337,1.1556113,-71.377727,-238.87507)"
       clip-path="url(#clipPath181-8)" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9);paint-order:fill markers stroke"
       d="m 72.907572,132.23981 0.313514,4.07981"
       id="path35-7"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-5);paint-order:fill markers stroke"
       d="m 76.926099,139.94821 3.035368,1.24454"
       id="path35-7-1"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-1);paint-order:fill markers stroke"
       d="m 87.535233,139.94638 -0.140128,3.28593"
       id="path35-7-0"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-16);paint-order:fill markers stroke"
       d="m 93.447344,137.82972 2.014673,-2.61142"
       id="path35-7-96"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#550000;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-0);paint-order:fill markers stroke"
       d="m 81.117505,135.75637 3.3756,-1.93095"
       id="path35-7-2"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#002e2e;stroke-width:0.785895;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-7);paint-order:fill markers stroke"
       d="m 82.272167,146.93618 -0.707181,1.92501"
       id="path35-7-6"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#000000;fill-opacity:0.972549;fill-rule:evenodd;stroke:#000000;stroke-width:1.4155;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-0-6);paint-order:fill markers stroke"
       d="m 80.928557,136.24066 5.927516,17.59103"
       id="path35-7-2-3"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#000000;fill-opacity:0.972549;fill-rule:evenodd;stroke:#000000;stroke-width:1.15265;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle-9-0-6-8);paint-order:fill markers stroke"
       d="M 136.27509,91.038238 122.51896,85.13419"
       id="path35-7-2-3-50"
       sodipodi:nodetypes="cc" />
    <path
       style="fill:#008080;fill-opacity:0.972549;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:1.00254;stroke-linecap:butt;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-start:url(#marker227);marker-end:url(#Stop);paint-order:fill markers stroke"
       d="m 82.976281,118.47623 13.602299,4.82732"
       id="path35-7-2-3-5"
       sodipodi:nodetypes="cc" />
    <g
       transform="matrix(0.77747678,0,0,0.77747678,90.734118,149.07577)"
       ns58:version="1.11.1"
       ns58:texconverter="pdflatex"
       ns58:pdfconverter="inkscape"
       ns58:text="$\\mathbf{u}$"
       ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
       ns58:scale="1.6424943957468967"
       ns58:alignment="middle center"
       ns58:inkscapeversion="1.4.2"
       ns58:jacobian_sqrt="0.579436"
       id="g225">
      <defs
         id="id-4ee86f0d-bc3c-4581-aadf-7996930d70ea" />
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-f5569139-3a6d-4661-8565-36c176759a34"
         transform="translate(-149.165,-130.281)">
        <g
           transform="translate(148.712,134.765)"
           id="g224">
          <path
             d="M 4.359375,-0.71875 V 0.0625 L 6.125,0 v -0.46875 c -0.609375,0 -0.6875,0 -0.6875,-0.390625 v -3.625 L 3.625,-4.40625 v 0.46875 c 0.609375,0 0.6875,0 0.6875,0.390625 v 1.90625 c 0,0.8125 -0.515625,1.34375 -1.234375,1.34375 -0.78125,0 -0.8125,-0.25 -0.8125,-0.796875 v -3.390625 l -1.8125,0.078125 v 0.46875 c 0.609375,0 0.6875,0 0.6875,0.390625 v 2.328125 c 0,1.0625 0.796875,1.28125 1.796875,1.28125 0.25,0 0.96875,0 1.421875,-0.78125 z m 0,0"
             id="id-192f29b4-9f2b-4cb6-8f72-1082341d0cb5" />
        </g>
      </g>
    </g>
    <g
       transform="matrix(0.84235494,0,0,0.84235494,89.624513,112.42774)"
       ns58:version="1.11.1"
       ns58:texconverter="pdflatex"
       ns58:pdfconverter="inkscape"
       ns58:text="$L$"
       ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
       ns58:scale="1.6424943957468967"
       ns58:alignment="middle center"
       ns58:inkscapeversion="1.4.2"
       ns58:jacobian_sqrt="0.579436"
       id="g227">
      <defs
         id="id-c06c0e0f-b6a9-406b-a1be-67048db7069a" />
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-55121ade-4086-4f63-9875-9b231a36d9b0"
         transform="translate(-149.103,-127.953)">
        <g
           transform="translate(148.712,134.765)"
           id="g226">
          <path
             d="M 3.734375,-6.03125 C 3.8125,-6.390625 3.84375,-6.5 4.78125,-6.5 c 0.296875,0 0.375,0 0.375,-0.1875 0,-0.125 -0.109375,-0.125 -0.15625,-0.125 -0.328125,0 -1.140625,0.03125 -1.46875,0.03125 -0.296875,0 -1.03125,-0.03125 -1.328125,-0.03125 -0.0625,0 -0.1875,0 -0.1875,0.203125 0,0.109375 0.09375,0.109375 0.28125,0.109375 0.015625,0 0.203125,0 0.375,0.015625 0.171875,0.03125 0.265625,0.03125 0.265625,0.171875 0,0.03125 0,0.0625 -0.03125,0.1875 L 1.5625,-0.78125 c -0.09375,0.390625 -0.109375,0.46875 -0.90625,0.46875 -0.171875,0 -0.265625,0 -0.265625,0.203125 C 0.390625,0 0.484375,0 0.65625,0 h 4.625 C 5.515625,0 5.515625,0 5.578125,-0.171875 L 6.375,-2.328125 c 0.03125,-0.109375 0.03125,-0.125 0.03125,-0.140625 0,-0.03125 -0.03125,-0.109375 -0.109375,-0.109375 -0.09375,0 -0.109375,0.0625 -0.171875,0.21875 -0.34375,0.90625 -0.78125,2.046875 -2.5,2.046875 H 2.6875 c -0.140625,0 -0.171875,0 -0.21875,0 -0.109375,-0.015625 -0.140625,-0.03125 -0.140625,-0.109375 0,-0.03125 0,-0.046875 0.046875,-0.21875 z m 0,0"
             id="id-be7987d1-295a-4536-b686-e5de29c88389" />
        </g>
      </g>
    </g>
    <g
       transform="matrix(0.69604788,0.00105675,-0.00105675,0.69604788,124.46646,76.574733)"
       ns58:version="1.11.1"
       ns58:texconverter="pdflatex"
       ns58:pdfconverter="inkscape"
       ns58:text="$\\mathbf{F_m}$"
       ns58:preamble="/home/bensabat/.config/inkscape/extensions/textext/default_packages.tex"
       ns58:scale="1.6424943957468967"
       ns58:alignment="middle center"
       ns58:inkscapeversion="1.4.2"
       ns58:jacobian_sqrt="0.579436"
       id="g236">
      <defs
         id="id-d4eab598-82c9-4dd7-900a-6485746f9c13" />
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-69034a1d-c836-45bc-808d-57cbea6c663f"
         transform="translate(-149.103,-127.984)">
        <g
           transform="translate(148.712,134.765)"
           id="g234">
          <path
             d="M 6.421875,-6.78125 H 0.390625 V -6.3125 H 1.46875 v 5.84375 H 0.390625 V 0 c 0.375,-0.03125 1.390625,-0.03125 1.828125,-0.03125 0.484375,0 1.5625,0 2.015625,0.03125 V -0.46875 H 2.875 v -2.6875 h 0.5 c 0.96875,0 1.046875,0.421875 1.046875,1.15625 h 0.46875 V -4.796875 H 4.421875 C 4.421875,-4.0625 4.34375,-3.625 3.375,-3.625 h -0.5 v -2.6875 h 1.40625 c 1.59375,0 1.828125,0.765625 1.984375,1.9375 h 0.46875 z m 0,0"
             id="id-6acd6b9b-93cc-4b0f-899a-8e9d41389feb" />
        </g>
      </g>
      <g
         fill="#000000"
         fill-opacity="1"
         id="id-cf94fed9-c7e5-40d7-834b-c3b6cec3f7b1"
         transform="translate(-149.103,-127.984)">
        <g
           transform="translate(155.921,136.259)"
           id="g235">
          <path
             d="m 6.75,-2.09375 c 0,-0.875 -0.578125,-1.046875 -1.203125,-1.046875 -0.65625,0 -1.09375,0.3125 -1.3125,0.65625 -0.171875,-0.609375 -0.78125,-0.65625 -1.15625,-0.65625 -0.828125,0 -1.234375,0.5 -1.375,0.734375 v -0.734375 l -1.25,0.0625 V -2.6875 c 0.40625,0 0.453125,0 0.453125,0.265625 v 2.03125 H 0.453125 V 0 c 0,0 0.5625,-0.03125 0.90625,-0.03125 C 1.6875,-0.03125 2.265625,0 2.265625,0 v -0.390625 h -0.46875 v -1.34375 c 0,-0.828125 0.75,-1.078125 1.140625,-1.078125 0.3125,0 0.453125,0.15625 0.453125,0.671875 v 1.75 H 2.921875 V 0 c 0,0 0.5625,-0.03125 0.90625,-0.03125 0.34375,0 0.90625,0.03125 0.90625,0.03125 v -0.390625 h -0.46875 v -1.34375 c 0,-0.828125 0.75,-1.078125 1.15625,-1.078125 0.3125,0 0.4375,0.15625 0.4375,0.671875 v 1.75 H 5.390625 V 0 C 5.40625,0 5.96875,-0.03125 6.296875,-0.03125 6.640625,-0.03125 7.203125,0 7.21875,0 V -0.390625 H 6.75 Z m 0,0"
             id="id-c6b34bc7-5c65-4524-8e78-4e69486596e8" />
        </g>
      </g>
    </g>
    <path
       d="M 60.349037,120.59789 48.313366,77.431557"
       style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
       id="path1-0"
       sodipodi:nodetypes="cc" />
    <path
       d="M 62.277314,70.689192 82.035036,105.77497"
       style="fill:#1a1a1a;fill-rule:evenodd;stroke:#1a1a1a;stroke-width:0.294635;stroke-linecap:round;stroke-linejoin:bevel;stroke-dasharray:none;stroke-dashoffset:0;paint-order:fill markers stroke"
       id="path1-03"
       sodipodi:nodetypes="cc" />
    <path
       style="opacity:1;fill:#800000;fill-opacity:0.972549;fill-rule:evenodd;stroke:#800000;stroke-width:0.745251;stroke-linecap:round;stroke-linejoin:round;stroke-dasharray:none;stroke-opacity:0.960784;marker-end:url(#ConcaveTriangle);paint-order:fill markers stroke"
       d="m 142.30215,93.491 -12.8098,-5.232214"
       id="path35" />
  </g>
</svg>
